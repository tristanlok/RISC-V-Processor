package riscV_pkg;
	import uvm_pkg::*;

	
endpackage
