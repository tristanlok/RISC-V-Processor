module control_unit (
	input [31:0]	instruction,
	
	output			reg_alu_mux,
	output			mem_read,
	output			mem_write,
	output [1:0]	alu_op,
	output			reg_write,
	output			data_reg_mux,
	output			branch_ctrl
);

assign 

endmodule
