 module riscv_top (
    input   logic       clk_in
);

    

endmodule
